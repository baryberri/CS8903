// Systolic Array's Size; 'N' means 'N x N' Systolic Array.
typedef 8 SystolicArraySize;
