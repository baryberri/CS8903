// Systolic Array's Size; 'N' means 'N x N' Systolic Array.
typedef 4 SystolicArraySize;

// Fixed-Point Numbers Quantization Factors
typedef 8 IntegerBits;
typedef 8 FractionBits;
