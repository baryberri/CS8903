typedef 4 SystolicArraySize;
