typedef Bit#(32) Data;
