import FixedPoint::*;

// Integer and Fraction Bits
typedef 8 IntegerBit;
typedef 8 FractionBit;


// Defined data type
typedef FixedPoint#(IntegerBit, FractionBit) FixedPointData;
