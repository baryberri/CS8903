module mkTestBench();

    // TODO: Fill in here

endmodule