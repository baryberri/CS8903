import Fifo::*;

import FP8::*;


interface FP8Adder;
    method Action putArgA(FP8 newArgA);
    method Action putArgB(FP8 newArgB);
    method ActionValue#(FP8) getResult();
endinterface

(* synthesize *)
module mkFP8Adder(FP8Adder);
    /*** Input and Output Fifos ***/
    Fifo#(1, FP8) argA <- mkBypassFifo();
    Fifo#(1, FP8) argB <- mkBypassFifo();

    Fifo#(1, FP8) result <- mkPipelineFifo();

    
    /*** Pipelining Fifos ***/
    Fifo#(1, FP8AdderOperands) decoded <- mkPipelineFifo();
    Fifo#(1, FP8AdderOperand) added <- mkPipelineFifo();
    Fifo#(1, FP8AdderOperand) shiftedBy2 <- mkPipelineFifo();
    Fifo#(1, FP8AdderOperand) shiftedBy1 <- mkPipelineFifo();


    /*** Rules ***/
    rule decode;
        // fetch
        let a = argA.first();
        let b = argB.first();

        argA.deq();
        argB.deq();

        // decode
        FP8AdderOperands operands = ?;

        operands.a.sign = a[7];
        operands.b.sign = b[7];

        operands.a.exponent = a[6:3];
        operands.b.exponent = b[6:3];

        if (operands.a.exponent == 0) begin
            // Denormal value
            operands.a.state = Normal;  // But we set this to Normal, because we manually set the exponent and mantissa correctly.
            operands.a.exponent = 1;
            operands.a.mantissa = {2'b00, a[2:0]};
        end else if (operands.a.exponent == '1) begin
            if (a[2:0] == 0) begin
                operands.a.state = Inf;
            end else begin
                operands.a.state = NaN;
            end
        end else begin
            // Normal value
            operands.a.state = Normal;
            operands.a.mantissa = {2'b01, a[2:0]};
        end

        if (operands.b.exponent == 0) begin
            operands.b.state = Normal;
            operands.b.exponent = 1;
            operands.b.mantissa = {2'b00, b[2:0]};
        end else if (operands.b.exponent == '1) begin
            if (b[2:0] == 0) begin
                operands.b.state = Inf;
            end else begin
                operands.b.state = NaN;
            end
        end else begin
            operands.b.state = Normal;
            operands.b.mantissa = {2'b01, b[2:0]};
        end

        // Match exponent
        if (operands.a.state == Normal && operands.b.state == Normal) begin
            if (operands.a.exponent >= operands.b.exponent) begin
                operands.b.mantissa = operands.b.mantissa >> (operands.a.exponent - operands.b.exponent);
                operands.b.exponent = operands.a.exponent;
            end else begin
                operands.a.mantissa = operands.a.mantissa >> (operands.b.exponent - operands.a.exponent);
                operands.a.exponent = operands.b.exponent;
            end
        end

        decoded.enq(operands);
    endrule

    rule addition;
        let operands = decoded.first();
        decoded.deq();
        
        FP8AdderOperand nextResult = ?;

        // Compute
        if (operands.a.state == Normal && operands.b.state == Normal) begin
            // Normal case
            nextResult.state = Normal;

            nextResult.exponent = operands.a.exponent;

            if (operands.a.sign == operands.b.sign) begin
                nextResult.sign = operands.a.sign;
                nextResult.mantissa = operands.a.mantissa + operands.b.mantissa;
            end else begin
                if (operands.a.mantissa > operands.b.mantissa) begin
                    nextResult.sign = operands.a.sign;
                    nextResult.mantissa = operands.a.mantissa - operands.b.mantissa;
                end else if (operands.a.mantissa < operands.b.mantissa) begin
                    nextResult.sign = operands.b.sign;
                    nextResult.mantissa = operands.b.mantissa - operands.a.mantissa;
                end else begin
                    nextResult.sign = 1'b0;
                    nextResult.mantissa = 0;
                end
            end
        end else begin
            // Special cases
            if (operands.a.state == NaN || operands.b.state == NaN) begin
                nextResult.state = NaN;
            end else if (operands.a.state == Inf && operands.b.state == Inf) begin
                if (operands.a.sign == operands.b.sign) begin
                    nextResult.sign = operands.a.sign;
                    nextResult.state = Inf;
                end else begin
                    nextResult.state = NaN;
                end
            end else if (operands.a.state == Inf) begin
                nextResult.sign = operands.a.sign;
                nextResult.state = Inf; 
            end else begin
                nextResult.sign = operands.b.sign;
                nextResult.state = Inf;
            end
        end

        added.enq(nextResult);
    endrule

    rule shiftBy2;
        let operand = added.first();
        added.deq();

        if (operand.state == Normal) begin
            // Make 1 be in [4:2] if it's in [1:0]
            if (operand.mantissa < (1 << 2)) begin
                if (operand.exponent <= 2) begin
                    operand.mantissa = operand.mantissa << (operand.exponent - 1);
                    operand.state = Denormal; 
                end else begin
                    operand.mantissa = operand.mantissa << 2;
                    operand.exponent = operand.exponent - 2;
                end
            end
        end

        shiftedBy2.enq(operand);
    endrule

    rule shiftBy1;
        let operand = shiftedBy2.first();
        shiftedBy2.deq();

        if (operand.state == Normal) begin
            // Make 1 be in [4:3] if it's in [2]
            if (operand.mantissa < (1 << 3)) begin
                if (operand.exponent <= 1) begin
                    // operand.exponent is <= 1 already: no need to shift mantissa anymore
                    operand.state = Denormal;
                end else begin
                    operand.mantissa = operand.mantissa << 1;
                    operand.exponent = operand.exponent - 1;
                end
            end
        end

        shiftedBy1.enq(operand);
    endrule

    rule putResult;
        let operand = shiftedBy1.first();
        shiftedBy1.deq();

        if (operand.state == Normal) begin
            // 1 is in [4:3]
            if (operand.mantissa[4] == 1'b1) begin
                operand.exponent = operand.exponent + 1;
                result.enq({operand.sign, operand.exponent, operand.mantissa[3:1]});
            end else begin
                result.enq({operand.sign, operand.exponent, operand.mantissa[2:0]});
            end
        end else if (operand.state == Denormal) begin
            operand.exponent = 0;
            result.enq({operand.sign, operand.exponent, operand.mantissa[2:0]});
        end else if (operand.state == Inf) begin
            operand.exponent = '1;
            operand.mantissa = 0;
            result.enq({operand.sign, operand.exponent, operand.mantissa[2:0]});
        end else begin
            // NaN
            operand.sign = 1'b0;
            operand.exponent = '1;
            operand.mantissa = 1;
            result.enq({operand.sign, operand.exponent, operand.mantissa[2:0]});
        end
    endrule


    /*** interfaces ***/
    method Action putArgA(FP8 newArgA);
        argA.enq(newArgA);
    endmethod

    method Action putArgB(FP8 newArgB);
        argB.enq(newArgB);
    endmethod

    method ActionValue#(FP8) getResult();
        result.deq();
        return result.first();
    endmethod
endmodule
