typedef 8 SystolicArraySize;

typedef Bit#(TLog#(SystolicArraySize)) PE_ID;
typedef Bit#(TAdd#(TLog#(SystolicArraySize), 1)) SystolicArrayID;
