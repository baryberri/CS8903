module mkFixedPointExamples();

    // TODO: Fill in here
    
endmodule
