typedef 16 SystolicArraySize;
