typedef Bit#(64) Data;
